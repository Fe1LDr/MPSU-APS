package filenames_pkg;

  parameter INSTR_INIT_FILE_NAME = "lab_13_ps2_vga_instr.mem";
  parameter  DATA_INIT_FILE_NAME = "lab_13_ps2ascii_data.mem";

endpackage